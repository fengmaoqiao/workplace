
--------------------------------------------------------------------------------
-- End of file
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--       ------------      Project : WILD Modem 802.11a2
--    ,' GoodLuck ,'      RCSfile: pilot_scr_pkg.vhd,v   
--   '-----------'     Author: DR \*
--
--  Revision: 1.1   
--  Date: 1999.12.31
--  State: Exp  
--  Locker:   
--------------------------------------------------------------------------------
--
-- Description : Package for pilot_scr.
--
--------------------------------------------------------------------------------
--
--  Source: ./git/COMMON/IPs/WILD/MODEM802_11a2/TX_TOP/pilot_scr/vhdl/rtl/pilot_scr_pkg.vhd,v  
--  Log: pilot_scr_pkg.vhd,v  
-- Revision 1.1  2003/03/13 15:02:28  Dr.A
-- Initial revision
--
--
--------------------------------------------------------------------------------


--------------------------------------------------------------------------------
-- Library
--------------------------------------------------------------------------------
library IEEE; 
use IEEE.STD_LOGIC_1164.ALL; 


--------------------------------------------------------------------------------
-- Package
--------------------------------------------------------------------------------
package pilot_scr_pkg is


--------------------------------------------------------------------------------
-- Components list declaration done by <fb> script.
--------------------------------------------------------------------------------
----------------------
-- File: pilot_scr.vhd
----------------------
  component pilot_scr
  port (
    --------------------------------------
    -- Clocks & Reset
    --------------------------------------
    reset_n           : in std_logic; -- asynchronous reset.
    clk               : in std_logic; -- Module clock.
    --------------------------------------
    -- Controls
    --------------------------------------
    enable_i          : in  std_logic; -- TX path enable.
    pilot_ready_i     : in  std_logic;
    init_pilot_scr_i  : in  std_logic;
    --------------------------------------
    -- Data
    --------------------------------------
    pilot_scr_o       : out std_logic  -- Data for the 4 pilot carriers.
    
  );

  end component;



 
end pilot_scr_pkg;

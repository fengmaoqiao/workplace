
--------------------------------------------------------------------------------
-- End of file
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--       ------------      Project : WILD Modem 802.11a2
--    ,' GoodLuck ,'      RCSfile: preamble_gen_pkg.vhd,v   
--   '-----------'     Author: DR \*
--
--  Revision: 1.2   
--  Date: 1999.12.31
--  State: Exp  
--  Locker:   
--------------------------------------------------------------------------------
--
-- Description : Package for preamble_gen.
--
--------------------------------------------------------------------------------
--
--  Source: ./git/COMMON/IPs/WILD/MODEM802_11a2/TX_TOP/preamble_gen/vhdl/rtl/preamble_gen_pkg.vhd,v  
--  Log: preamble_gen_pkg.vhd,v  
-- Revision 1.2  2003/10/13 09:42:55  Dr.B
-- Corrected long_seq_re(23): was coded -86 is now -82.
--
-- Revision 1.1  2003/03/13 15:04:58  Dr.A
-- Initial revision
--
--
--------------------------------------------------------------------------------


--------------------------------------------------------------------------------
-- Library
--------------------------------------------------------------------------------
library IEEE; 
use IEEE.STD_LOGIC_1164.ALL; 


--------------------------------------------------------------------------------
-- Package
--------------------------------------------------------------------------------
package preamble_gen_pkg is

  ------------------------------------------------------------------------------
  -- Types
  ------------------------------------------------------------------------------
  type integer_ar_16 is array (0 to 15) of std_logic_vector(9 downto 0);
  type integer_ar_32 is array (0 to 31) of std_logic_vector(9 downto 0);

  ------------------------------------------------------------------------------
  -- Constants
  ------------------------------------------------------------------------------
  
  -- ROMS for short and long preamble symbols i and q values.
  
  -- Short training sequence
  constant short_seq_re : integer_ar_16 := (
    "0001000011", -- 67,
    "1100111111", -- -193, 
    "1111101100", -- -20, 
    "0011010000", -- 208, 
    "0010000110", -- 134, 
    "0011010000", -- 208, 
    "1111101100", -- -20,
    "1100111111", -- -193, 
    "0001000011", -- 67, 
    "0000000011", -- 3, 
    "1110001110", -- -114, 
    "1111101110", -- -18, 
    "0000000000", -- 0, 
    "1111101110", -- -18,
    "1110001110", -- -114, 
    "0000000011"  -- 3, 
    );

  constant short_seq_im : integer_ar_16 := (
    "0001000011", -- 67, 
    "0000000011", -- 3, 
    "1110001110", -- -114, 
    "1111101110", -- -18, 
    "0000000000", -- 0, 
    "1111101110", -- -18, 
    "1110001110", -- -114, 
    "0000000011", -- 3, 
    "0001000011", -- 67, 
    "1100111111", -- -193, 
    "1111101100", -- -20, 
    "0011010000", -- 208, 
    "0010000110", -- 134, 
    "0011010000", -- 208, 
    "1111101100", -- -20,
    "1100111111" -- -193
    );

  -- Long training sequence
  constant long_seq_re : integer_ar_32 := (
    "0011100100", -- 228, 
    "1111111001", -- -7, 
    "0000111010", -- 58, 
    "0010001101", -- 141, 
    "0000011111", -- 31, 
    "0001010111", -- 87, 
    "1101011000", -- -168, 
    "1111001000", -- -56,
    "0010001110", -- 142, 
    "0001001110", -- 78, 
    "0000000001", -- 1, 
    "1100111001", -- -199, 
    "0000100100", -- 36, 
    "0001010101", -- 85, 
    "1111011111", -- -33, 
    "0010101110", -- 174,
    "0001011011", -- 91, 
    "0000110110", -- 54, 
    "1110101101", -- -83, 
    "1101000001", -- -191, 
    "0001111000", -- 120, 
    "0001100101", -- 101, 
    "1110101000", -- -88,
    "1110101110", -- -82, 
    "1111001101", -- -51, 
    "1101001111", -- -177, 
    "1101000111", -- -185, 
    "0001101101", -- 109, 
    "1111111100", -- -4, 
    "1101111010", -- -134,
    "0010000110", -- 134, 
    "0000010010" -- 18, 
    );

  constant long_seq_im : integer_ar_32 := (
    "0000000000",  -- 0, 
    "1101010001", -- -175, 
    "1101011110", -- -162, 
    "0001111001", -- 121, 
    "0000101001", -- 41, 
    "1110000000", -- -128, 
    "1110110000", -- -80,
    "1101100101", -- -155, 
    "1111011010", -- -38, 
    "0000000110", -- 6, 
    "1101011001", -- -167, 
    "1110111011", -- -69, 
    "1110101011", -- -85, 
    "1111101010", -- -22,
    "0011101010", -- 234, 
    "1111111010", -- -6, 
    "1110100101", -- -91, 
    "0010001111", -- 143, 
    "0000111001", -- 57, 
    "0001011111", -- 95, 
    "0010000110", -- 134,
    "0000010101", -- 21,
    "0001110110", -- 118, 
    "1111100000", -- -32, 
    "1100100100", -- -220, 
    "1111101000", -- -24, 
    "1111100010", -- -30, 
    "1110010100", -- -108, 
    "0001001110", -- 78, 
    "0010101000", -- 168, 
    "0010011010", -- 154, 
    "0010001110"  -- 142, 
    );

--------------------------------------------------------------------------------
-- Components list declaration done by <fb> script.
--------------------------------------------------------------------------------
----------------------
-- File: preamble_gen.vhd
----------------------
  component preamble_gen
  port (
    --------------------------------------
    -- Clocks & Reset
    --------------------------------------
    clk             : in  std_logic; -- Module clock
    reset_n         : in  std_logic; -- Asynchronous reset
    --------------------------------------
    -- Controls
    --------------------------------------
    enable_i        : in  std_logic; -- TX path enable.
    data_ready_i    : in  std_logic; -- '1' when next block ready to accept data
    add_short_pre_i : in  std_logic_vector(1 downto 0); -- pre-preamble value.
    --
    end_preamble_o  : out std_logic; -- High at the end of the preamble.
    --------------------------------------
    -- Data
    --------------------------------------
    i_out           : out std_logic_vector(9 downto 0); -- I preamble data.
    q_out           : out std_logic_vector(9 downto 0)  -- Q preamble data.
  );

  end component;



 
end preamble_gen_pkg;

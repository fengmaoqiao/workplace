
--------------------------------------------------------------------------------
-- End of file
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--       ------------      Project : bit_ser_adder
--    ,' GoodLuck ,'      RCSfile: fa.vhd,v  
--   '-----------'     Author: DR \*
--
--  Revision: 1.1  
--  Date: 1999.12.31
--  State: Exp  
--  Locker:   
--------------------------------------------------------------------------------
--
-- Description : Full adder
--
--
--------------------------------------------------------------------------------
--
--  Source: ./git/COMMON/IPs/NLWARE/DSP/bit_ser_adder/vhdl/rtl/fa.vhd,v  
--  Log: fa.vhd,v  
-- Revision 1.1  2003/04/18 07:07:54  rrich
-- Initial revision
--
--
--
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Library
--------------------------------------------------------------------------------
library IEEE; 
use IEEE.STD_LOGIC_1164.ALL;

--library bit_ser_adder_rtl;
library work;
--use bit_ser_adder_rtl.bit_ser_adder_pkg.all;
use work.bit_ser_adder_pkg.all;

--------------------------------------------------------------------------------
-- Entity
--------------------------------------------------------------------------------
entity fa is
  
  port (
    x     : in  std_logic;
    y     : in  std_logic;
    c_in  : in  std_logic;
    s     : out std_logic;
    c_out : out std_logic);

end fa;

--------------------------------------------------------------------------------
-- Architecture
--------------------------------------------------------------------------------
architecture rtl of fa is

  ------------------------------------------------------------------------------
  -- Signals
  ------------------------------------------------------------------------------
  signal c_0, c_1, s_0 : std_logic;
  
begin  -- rtl

  ha_0 : ha
    port map (
      x => x,
      y => y,
      c => c_0,
      s => s_0);
     
  ha_1 : ha
    port map (
      x => s_0,
      y => c_in,
      c => c_1,
      s => s);

  c_out <= c_0 or c_1;

end rtl;




--------------------------------------------------------------------------------
-- End of file
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--       ------------      Project : WiLDBuP2
--    ,' GoodLuck ,'      RCSfile: mem2_seq_pkg.vhd,v  
--   '-----------'     Author: DR \*
--
--  Revision: 1.5  
--  Date: 1999.12.31
--  State: Exp  
--  Locker:   
--------------------------------------------------------------------------------
--
-- Description : Package for mem2_seq.
--
--------------------------------------------------------------------------------
--
--  Source: ./git/COMMON/IPs/WILD/WILDBuP2/mem2_seq/vhdl/rtl/mem2_seq_pkg.vhd,v  
--  Log: mem2_seq_pkg.vhd,v  
-- Revision 1.5  2005/05/31 15:51:23  Dr.A
-- #BugId:938#
-- Removed unused signals
--
-- Revision 1.4  2005/02/09 17:54:06  Dr.A
-- #BugId:974#
-- Reset_bufempty sent on RX write access
--
-- Revision 1.3  2004/04/14 16:06:08  Dr.A
-- Removed unused signal last_word_size.
--
-- Revision 1.2  2004/01/26 08:50:22  Dr.F
-- added ready_load.
--
-- Revision 1.1  2003/11/19 16:27:34  Dr.F
-- Initial revision
--
--
--------------------------------------------------------------------------------


--------------------------------------------------------------------------------
-- Library
--------------------------------------------------------------------------------
library IEEE; 
    use IEEE.STD_LOGIC_1164.ALL; 


--------------------------------------------------------------------------------
-- Package
--------------------------------------------------------------------------------
package mem2_seq_pkg is


--------------------------------------------------------------------------------
-- Components list declaration done by <fb> script.
--------------------------------------------------------------------------------

 
end mem2_seq_pkg;
